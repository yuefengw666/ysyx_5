module ysyx_22040237_ifu(
  //input clk,
  //input rst,
  input [31:0] inst_i,
  output [31:0] inst_o
);

assign inst_o = inst_i;

endmodule
